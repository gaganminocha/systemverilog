`timescale 1ns/100ps
`include full_adder.sv

module full_adder_tb;
	reg 



endmodule
